module or_gate(a,b,z);
input a,b;
output z;

assign z=a|b;

endmodule